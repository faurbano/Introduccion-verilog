//-- Prueba FPGA IceZum Alhambra
module leds(output wire LED0,
            output wire LED1);

//-- Asignación LEDS
assign LED0 = 1'b1;
assign LED1 = 1'b1;

endmodule
